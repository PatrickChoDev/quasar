`include "./fp.vh"
